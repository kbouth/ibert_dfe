
// file: ibert_test.v
//////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2012.3
//  \   \         Application : IBERT 7Series 
//  /   /         Filename : example_ibert_ultrascale_gth_0
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module ibert_test
// Generated by Xilinx IBERT_7S 
//////////////////////////////////////////////////////////////////////////////

`define C_NUM_GTH_QUADS 2
`define C_GTH_REFCLKS_USED 1
module ibert_test
(
  // GT top level ports
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txn_o,
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txp_o,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]    	gth_rxn_i,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]   	gth_rxp_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0n_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1n_i,
    output                                sys_clk_debug, 
  output                                sys_clk_buf, 
  output                                ref_clk_buf
);

  //
  // Ibert refclk internal signals
  //
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk1_i;        	
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk11_i; 
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk1_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_1_i;
  wire                        gth_sysclk_i;

  wire      clk; 
  wire                                   sys_clk;

   top system(
    .pl_clk0(sys_clk)
   );
   
  //
  // Refclk IBUFDS instantiations
  //
    IBUFDS_GTE4 u_buf_gth_q1_clk0
      (
        .O            (gth_refclk0_i[0]),
        .ODIV2        (gth_odiv2_0_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[0]),
        .IB           (gth_refclk0n_i[0])
      );

    IBUFDS_GTE4 u_buf_gth_q1_clk1
      (
        .O            (gth_refclk1_i[0]),
        .ODIV2        (gth_odiv2_1_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[0]),
        .IB           (gth_refclk1n_i[0])
      );
      
    BUFG_GT #(
       .SIM_DEVICE("ULTRASCALE_PLUS")  // ULTRASCALE, ULTRASCALE_PLUS
    )
    BUFG_GT_inst (
       .O(ref_clk_buf),             // 1-bit output: Buffer
       .CE(1'b1),           // 1-bit input: Buffer enable
       .CEMASK(1'b0),   // 1-bit input: CE Mask
       .CLR(1'b0),         // 1-bit input: Asynchronous clear
       .CLRMASK(1'b0), // 1-bit input: CLR Mask
       .DIV(3'b000),         // 3-bit input: Dynamic divide Value
       .I(gth_odiv2_1_i[0])              // 1-bit input: Buffer
    );
      
     sys_clk sys_clk0(
        .clk_in1(sys_clk),
        .clk_out1(clk)
    );
  //
  // Refclk connection from each IBUFDS to respective quads depending on the source selected in gui
  //
  assign gth_qrefclk0_i[0] = gth_refclk0_i[0];
  assign gth_qrefclk1_i[0] = gth_refclk1_i[0];
  assign gth_qnorthrefclk0_i[0] = 1'b0;
  assign gth_qnorthrefclk1_i[0] = 1'b0;
  assign gth_qsouthrefclk0_i[0] = 1'b0;
  assign gth_qsouthrefclk1_i[0] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[0] = gth_refclk0_i[0];
  assign gth_qrefclk10_i[0] = gth_refclk1_i[0];
  assign gth_qrefclk01_i[0] = gth_refclk0_i[0];
  assign gth_qrefclk11_i[0] = gth_refclk1_i[0];
  assign gth_qnorthrefclk00_i[0] = 1'b0;
  assign gth_qnorthrefclk10_i[0] = 1'b0;
  assign gth_qnorthrefclk01_i[0] = 1'b0;
  assign gth_qnorthrefclk11_i[0] = 1'b0;  
  assign gth_qsouthrefclk00_i[0] = 1'b0;
  assign gth_qsouthrefclk10_i[0] = 1'b0;  
  assign gth_qsouthrefclk01_i[0] = 1'b0;
  assign gth_qsouthrefclk11_i[0] = 1'b0; 
  assign sys_clk_debug = clk; 
  assign sys_clk_buf = clk;
  assign gth_qrefclk0_i[1] = 1'b0;
  assign gth_qrefclk1_i[1] = 1'b0;
  assign gth_qnorthrefclk0_i[1] = gth_refclk0_i[0];
  assign gth_qnorthrefclk1_i[1] = 1'b0;
  assign gth_qsouthrefclk0_i[1] = 1'b0;
  assign gth_qsouthrefclk1_i[1] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[1] = 1'b0;
  assign gth_qrefclk10_i[1] = 1'b0;
  assign gth_qrefclk01_i[1] = 1'b0;
  assign gth_qrefclk11_i[1] = 1'b0;
  assign gth_qnorthrefclk00_i[1] = gth_refclk0_i[0];
  assign gth_qnorthrefclk10_i[1] = 1'b0;
  assign gth_qnorthrefclk01_i[1] = gth_refclk0_i[0];
  assign gth_qnorthrefclk11_i[1] = 1'b0;
  assign gth_qsouthrefclk00_i[1] = 1'b0;
  assign gth_qsouthrefclk10_i[1] = 1'b0;
  assign gth_qsouthrefclk01_i[1] = 1'b0;
  assign gth_qsouthrefclk11_i[1] = 1'b0;
  //
  // Sysclock connection
  //


  //
  // IBERT core instantiation
  //
  ibert u_ibert_gth_core
    (
      .txn_o(gth_txn_o),
      .txp_o(gth_txp_o),
      .rxn_i(gth_rxn_i),
      .rxp_i(gth_rxp_i),
      .clk(clk),
      .gtrefclk0_i(gth_qrefclk0_i),
      .gtrefclk1_i(gth_qrefclk1_i),
      .gtnorthrefclk0_i(gth_qnorthrefclk0_i),
      .gtnorthrefclk1_i(gth_qnorthrefclk1_i),
      .gtsouthrefclk0_i(gth_qsouthrefclk0_i),
      .gtsouthrefclk1_i(gth_qsouthrefclk1_i),
      .gtrefclk00_i(gth_qrefclk00_i),
      .gtrefclk10_i(gth_qrefclk10_i),
      .gtrefclk01_i(gth_qrefclk01_i),
      .gtrefclk11_i(gth_qrefclk11_i),
      .gtnorthrefclk00_i(gth_qnorthrefclk00_i),
      .gtnorthrefclk10_i(gth_qnorthrefclk10_i),
      .gtnorthrefclk01_i(gth_qnorthrefclk01_i),
      .gtnorthrefclk11_i(gth_qnorthrefclk11_i),
      .gtsouthrefclk00_i(gth_qsouthrefclk00_i),
      .gtsouthrefclk10_i(gth_qsouthrefclk10_i),
      .gtsouthrefclk01_i(gth_qsouthrefclk01_i),
      .gtsouthrefclk11_i(gth_qsouthrefclk11_i)
    );

endmodule

